
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:05:18 11/16/2017 
// Design Name: 
// Module Name:    digits_to_segments 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module digits_to_segments(
								clk,
								thousands,
								hundreds,
								tens,
								ones,
								thousands_segs,
								hundreds_segs,
								tens_segs,
								ones_segs
    );
	/////////////////////////////////////////////////////////////////////////////////
	//Inputs/Outputs
	/////////////////////////////////////////////////////////////////////////////////
	input clk;
   input [3:0] thousands;
   input [3:0] hundreds;
   input [3:0] tens;
   input [3:0] ones;
   output [7:0] thousands_segs;
   output [7:0] hundreds_segs;
   output [7:0] tens_segs;
   output [7:0] ones_segs;
	
	/////////////////////////////////////////////////////////////////////////////////
	//Wire/Reg Declarations
	/////////////////////////////////////////////////////////////////////////////////
	
	/////////////////////////////////////////////////////////////////////////////////
	//Constants
	/////////////////////////////////////////////////////////////////////////////////
	
	/////////////////////////////////////////////////////////////////////////////////
	//Sequential Logic
	/////////////////////////////////////////////////////////////////////////////////
	
	/////////////////////////////////////////////////////////////////////////////////
	//Module Instantiations
	/////////////////////////////////////////////////////////////////////////////////
	convert_to_segments a(thousands, thousands_segs);
	convert_to_segments b(hundreds, hundreds_segs);
	convert_to_segments c(tens, tens_segs);
	convert_to_segments d(ones, ones_segs);
endmodule
